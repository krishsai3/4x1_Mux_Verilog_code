module mux_4_1 ( a, b, c, d, s0, s1, out);

input wire a, b, c, d;
input wire s0, s1;
output reg out;

always @ (a or b or c or d or s0, s1)
begin

case (s0 | s1)
2'b00 : out <= a;
2'b01 : out <= b;
2'b10 : out <= c;
2'b11 : out <= d;
endcase

end

endmodule

//testbench
module mux_4_1_tb;
    wire  out;
    reg  a;
    reg  b;
    reg  c;
    reg  d;
    reg s0, s1;

mux_4_1 mux(.a(a),.b(b),.c(c),.d(d),.s0(s0),.s1(s1),out(out));

initial
    begin
     a=1'b0; 
     b=1'b0; 
     c=1'b0; 
     d=1'b0;
     s0=1'b0; 
     s1=1'b0;
     #500 $finish;
    end
always #40 a=~a;
always #20 b=~b;
always #10 c=~c;
always #5 d=~d;
always #80 s0=~s0;
always #160 s1=~s1;
    
always @(a or b or c or d or s0 or s1)
$monitor("At time =%t, Output%d",$time,out);

endmodule